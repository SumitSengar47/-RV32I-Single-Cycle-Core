`timescale 1ns/1ps

// This is a self-checking testbench for the extend.v module.
// It verifies that the immediate generator correctly extracts and sign-extends
// values for all supported RISC-V immediate formats.

module extend_tb;

    // --- DUT Signals ---
    reg  [31:0] instr;     // The 32-bit instruction to be decoded.
    reg  [2:0]  imm_src;   // The 3-bit control signal selecting the format.
    wire [31:0] imm_ext;   // The 32-bit immediate value generated by the DUT.

    // --- Instantiate the DUT (Device Under Test) ---
    extend dut (
        .instr(instr),
        .imm_src(imm_src),
        .imm_ext(imm_ext)
    );

    // --- Local Parameters for Control Signal ---
    // These codes must match the ones used in the main_decoder.
    localparam IMM_I = 3'd0; // I-type
    localparam IMM_S = 3'd1; // S-type
    localparam IMM_B = 3'd2; // B-type
    localparam IMM_U = 3'd3; // U-type
    localparam IMM_J = 3'd4; // J-type
    localparam IMM_R = 3'd5; // R-type (no immediate)

    // --- Verification Infrastructure ---
    integer total = 0;
    integer passed = 0;

    // --- Helper Task for Test Execution ---
    // This task applies a test vector, computes the expected result locally,
    // and compares it against the DUT's output.
    task run_case;
        input [31:0] t_instr;
        input [2:0]  t_imm_src;
        input [80:1] desc;
        reg   [31:0] expected;
        begin
            // Apply inputs to the DUT.
            instr   = t_instr;
            imm_src = t_imm_src;
            #2; // Allow a small delay for the combinational logic to settle.

            // This "golden model" calculates the expected result using the same
            // logic as the DUT, providing a reliable reference for comparison.
            case (t_imm_src)
                IMM_I: expected = {{20{instr[31]}}, instr[31:20]};
                IMM_S: expected = {{20{instr[31]}}, instr[31:25], instr[11:7]};
                IMM_B: expected = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
                IMM_U: expected = {instr[31:12], 12'b0};
                IMM_J: expected = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
                IMM_R: expected = 32'h00000000;
                default: expected = 32'h00000000;
            endcase

            // Compare the DUT's output with the expected value and report the result.
            total = total + 1;
            if (imm_ext === expected) begin
                passed = passed + 1;
                $display("%0t | PASS | %s | imm_src=%0d instr=0x%h -> imm_ext=0x%h",
                         $time, desc, t_imm_src, instr, imm_ext);
            end else begin
                $display("%0t | FAIL | %s | imm_src=%0d instr=0x%h -> got=0x%h expected=0x%h",
                         $time, desc, t_imm_src, instr, imm_ext, expected);
            end
            #1;
        end
    endtask

    // --- Test Sequence ---
    initial begin
        // Enable waveform dumping for visual debugging.
        $dumpfile("extend_tb.vcd");
        $dumpvars(0, extend_tb);

        // --- Test Vectors ---
        // Each vector is a full 32-bit instruction word, constructed by concatenating
        // the required fields according to the RISC-V specification.

        // Test I-type with a negative immediate (-4).
        instr = { 12'hFFC, 5'd9, 3'b010, 5'd6, 7'b0000011 };
        run_case(instr, IMM_I, "I-type lw (imm=-4)");

        // Test I-type with a positive immediate (8).
        instr = { 12'h008, 5'd1, 3'b000, 5'd2, 7'b0010011 };
        run_case(instr, IMM_I, "I-type addi (imm=8)");

        // Test S-type with a positive immediate (8).
        instr = { 7'b0000000, 5'd6, 5'd9, 3'b010, 5'b01000, 7'b0100011 };
        run_case(instr, IMM_S, "S-type sw (imm=8)");

        // Test B-type with a negative offset (-4).
        instr = { 1'b1, 6'b111111, 5'd4, 5'd4, 3'b000, 4'b1100, 1'b1, 7'b1100011 };
        run_case(instr, IMM_B, "B-type beq (offset = -4)");

        // Test U-type for LUI.
        instr = { 20'h12345, 5'd5, 7'b0110111 };
        run_case(instr, IMM_U, "U-type LUI (imm=0x12345<<12)");

        // Test J-type for JAL.
        instr = { 1'b0, 10'd1, 1'b0, 8'h01, 5'd1, 7'b1101111 };
        run_case(instr, IMM_J, "J-type JAL (small +offset)");

        // Test R-type (should produce a zero immediate).
        instr = 32'h0062E233; // An example R-type instruction.
        run_case(instr, IMM_R, "R-type (no immediate)");

        // --- Final Summary ---
        #5;
        $display("==== SUMMARY: %0d / %0d passed ====", passed, total);
        if (passed != total) $display("Some tests failed - inspect messages or extend_tb.vcd");
        else $display("All tests passed.");
        $finish;
    end

    // Optional monitor for continuous signal tracking.
    initial begin
        $monitor("t=%0t instr=0x%08h imm_src=%0d imm_ext=0x%08h", $time, instr, imm_src, imm_ext);
    end

endmodule
