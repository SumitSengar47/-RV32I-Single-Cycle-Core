// extend.v
// Immediate extender for a RISC-V processor.

// This module decodes the various immediate formats from the raw instruction bits.
// The `imm_src` input signal selects which format to extract and generate.

module extend (
    // --- Ports ---
    input  wire [31:0] instr,      // The full 32-bit instruction word.
    input  wire [2:0]  imm_src,    // A 3-bit control signal that selects the format.
    output reg  [31:0] imm_ext     // The final 32-bit sign-extended immediate value.
);

    // --- Local Parameters for Control Signal ---
    // These codes must match the ones generated by the main_decoder.
    localparam IMM_I = 3'd0; // I-type (e.g., ADDI, LW)
    localparam IMM_S = 3'd1; // S-type (e.g., SW)
    localparam IMM_B = 3'd2; // B-type (e.g., BEQ)
    localparam IMM_U = 3'd3; // U-type (e.g., LUI)
    localparam IMM_J = 3'd4; // J-type (e.g., JAL)
    localparam IMM_R = 3'd5; // R-type (no immediate)

    // --- Combinational Logic for Immediate Generation ---
    // This block is always active and will update the output whenever an input changes.
    always @(*) begin
        // The case statement selects the correct logic based on the control signal.
        case (imm_src)
            // I-type: sign-extend the 12-bit immediate from instr[31:20].
            IMM_I: imm_ext = {{20{instr[31]}}, instr[31:20]};

            // S-type: reconstruct and sign-extend the 12-bit immediate from two fields.
            IMM_S: imm_ext = {{20{instr[31]}}, instr[31:25], instr[11:7]};

            // B-type: reconstruct and sign-extend the 13-bit immediate for branches.
            IMM_B: imm_ext = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};

            // U-type: place the 20-bit immediate in the upper bits, zeroing the lower 12.
            IMM_U: imm_ext = {instr[31:12], 12'b0};

            // J-type: reconstruct and sign-extend the 21-bit immediate for jumps.
            IMM_J: imm_ext = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};

            // R-type or unused: return zero as there is no immediate.
            IMM_R: imm_ext = 32'h0000_0000;

            // A safe default to prevent latches.
            default: imm_ext = 32'h0000_0000;
        endcase
    end

endmodule

