// alu.v
// Combinational ALU for a RISC-V RV32I processor.
// - Implements arithmetic, logical, and shift operations.
// - Uses a robust, three-stage structure to prevent simulation hazards.

module alu (
    input  wire [31:0] src_a,         // ALU input A (from register file or PC)
    input  wire [31:0] src_b,         // ALU input B (from register file or immediate)
    input  wire [3:0]  alu_control,   // Operation select from the control unit
    output reg  [31:0] alu_result,    // The 32-bit result of the operation
    output wire        zero,          // Flag: set to 1 if alu_result is all zeros
    output wire        carry,         // Flag: carry-out from addition/subtraction
    output wire        overflow,      // Flag: signed overflow from addition/subtraction
    output wire        negative       // Flag: the most significant bit of alu_result
);

    // -------------------------------------------------------------------------
    // ALU Control Codes
    // -------------------------------------------------------------------------
    // These local parameters define the 4-bit codes for each ALU operation.
    // They must match the codes generated by the alu_decoder module.
    localparam ALU_ADD   = 4'b0000; // Addition (for ADD, ADDI)
    localparam ALU_SUB   = 4'b0001; // Subtraction (for SUB, and all branches)
    localparam ALU_AND   = 4'b0010; // Bitwise AND
    localparam ALU_OR    = 4'b0011; // Bitwise OR
    localparam ALU_XOR   = 4'b0100; // Bitwise XOR
    localparam ALU_SLT   = 4'b0101; // Set Less Than (signed)
    localparam ALU_SLTU  = 4'b0110; // Set Less Than (unsigned)
    localparam ALU_SLL   = 4'b0111; // Shift Left Logical
    localparam ALU_SRL   = 4'b1000; // Shift Right Logical
    localparam ALU_SRA   = 4'b1001; // Shift Right Arithmetic
    localparam ALU_LUI   = 4'b1010; // Load Upper Immediate (passthrough)
    localparam ALU_AUIPC = 4'b1011; // Add Upper Immediate to PC (uses adder)

    // -------------------------------------------------------------------------
    // Stage 1: Parallel Calculation Units
    // -------------------------------------------------------------------------
    // All possible results are calculated here in parallel *before* selection.
    // This robust design pattern prevents the combinatorial feedback loops
    // that caused X-propagation issues in previous versions.

    // An internal wire to determine if the current operation is a subtraction.
    // This simplifies the adder/subtractor logic below.
    wire is_sub = (alu_control == ALU_SUB);

    // A single, 33-bit wide adder/subtractor unit.
    // For subtraction (A-B), we compute A + (~B) + 1 using two's complement.
    // The 33rd bit (sum_wide[32]) correctly captures the carry-out.
    wire [32:0] sum_wide = {1'b0, src_a} + (is_sub ? {1'b0, ~src_b} : {1'b0, src_b}) + (is_sub ? 1'b1 : 1'b0);
    wire [31:0] add_sub_result = sum_wide[31:0];

    // The results for all logical, shift, and comparison operations are also calculated in parallel.
    wire [31:0] and_result  = src_a & src_b;
    wire [31:0] or_result   = src_a | src_b;
    wire [31:0] xor_result  = src_a ^ src_b;
    wire [31:0] slt_result  = ($signed(src_a) < $signed(src_b)) ? 32'd1 : 32'd0;
    wire [31:0] sltu_result = (src_a < src_b) ? 32'd1 : 32'd0;
    wire [31:0] sll_result  = src_a << src_b[4:0];
    wire [31:0] srl_result  = src_a >> src_b[4:0];
    wire [31:0] sra_result  = $signed(src_a) >>> src_b[4:0]; // Use Verilog's built-in signed shift

    // -------------------------------------------------------------------------
    // Stage 2: Final Result Multiplexer
    // -------------------------------------------------------------------------
    // This 'always' block acts as a pure multiplexer. It selects one of the
    // pre-calculated results from Stage 1 based on the alu_control signal.
    // This structure is guaranteed to prevent inferred latches.
    always @(*) begin
        case (alu_control)
            ALU_ADD, ALU_SUB, ALU_AUIPC: alu_result = add_sub_result;
            ALU_AND:  alu_result = and_result;
            ALU_OR:   alu_result = or_result;
            ALU_XOR:  alu_result = xor_result;
            ALU_SLT:  alu_result = slt_result;
            ALU_SLTU: alu_result = sltu_result;
            ALU_SLL:  alu_result = sll_result;
            ALU_SRL:  alu_result = srl_result;
            ALU_SRA:  alu_result = sra_result;
            ALU_LUI:  alu_result = src_b;         // For LUI, the ALU just passes the immediate value through.
            default:  alu_result = 32'hDEADBEEF; // A known garbage value helps spot errors during debug.
        endcase
    end

    // -------------------------------------------------------------------------
    // Stage 3: Flag Generation
    // -------------------------------------------------------------------------
    // All flags are generated from the final, stable alu_result and the original inputs.
    // This structure is guaranteed to be free of combinatorial loops.

    // The 'zero' flag is true if all 32 bits of the result are zero.
    assign zero     = (alu_result == 32'h0);
  
    // The 'negative' flag is simply the most significant bit (MSB) of the result.
    assign negative = alu_result[31];

    // *** BUG FIX HERE ***
    // The 'carry' flag is ONLY meaningful for add/sub operations.
    // It is now explicitly set to 0 for all other operations to prevent incorrect flag values.
    // For subtraction (A-B), a carry-out of 1 means *no borrow* (i.e., A >= B).
    assign carry = ((alu_control == ALU_ADD) || (alu_control == ALU_SUB) || (alu_control == ALU_AUIPC)) ? sum_wide[32] : 1'b0;

    // Signed overflow logic is only meaningful for add/sub operations.
    // It occurs if the sign of the result is different from the sign of the inputs
    // (when the inputs have the same sign).
    wire add_overflow = (~src_a[31] & ~src_b[31] &  add_sub_result[31]) |
                        ( src_a[31] &  src_b[31] & ~add_sub_result[31]);
    wire sub_overflow = (~src_a[31] &  src_b[31] &  add_sub_result[31]) |
                        ( src_a[31] & ~src_b[31] & ~add_sub_result[31]);

    // Select the correct overflow flag based on the current operation.
    assign overflow = ((alu_control == ALU_ADD) || (alu_control == ALU_AUIPC)) ? add_overflow :
                      (alu_control == ALU_SUB) ? sub_overflow :
                      1'b0; // Overflow is not defined for logical/shift ops.

endmodule

